`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:20:11 02/15/2018 
// Design Name: 
// Module Name:    Bitwise 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Bitwise(a, b, x);
	input wire [7:0] a;
	input wire [7:0] b;
	output wire [7:0] x;
	
	 

endmodule
