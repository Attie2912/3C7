`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:14:51 02/06/2018 
// Design Name: 
// Module Name:    BarrelShift 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BarrelShift(
	input wire [31:0] a,
	input wire [4:0] amt,
	output reg [31:0] y,
	input wire direction
    );

always @*
 begin
	 if(direction == 1) // left 
		case(amt)
			5'b00000: y = a;
			5'o1: y = {a[0], a[31:1]};
			5'o2: y = {a[1:0], a[31:2]};
			5'o3: y = {a[2:0], a[31:3]};
			5'o4: y = {a[3:0], a[31:4]};
			5'o5: y = {a[4:0], a[31:5]};
			5'o6: y = {a[5:0], a[31:6]};
			5'o7: y = {a[6:0], a[31:7]};
			5'o10: y = {a[7:0], a[31:8]};
			5'o11: y = {a[8:0], a[31:9]};
			5'o12: y = {a[9:0], a[31:10]};
			5'o13: y = {a[10:0], a[31:11]};
			5'o14: y = {a[11:0], a[31:12]};
			5'o15: y = {a[12:0], a[31:13]};//13
			5'o16: y = {a[13:0], a[31:14]};
			5'o17: y = {a[14:0], a[31:15]};
			5'o20: y = {a[15:0], a[31:16]};
			5'o21: y = {a[16:0], a[31:17]};
			5'o22: y = {a[17:0], a[31:18]};
			5'o23: y = {a[18:0], a[31:19]};
			5'o24: y = {a[19:0], a[31:20]};
			5'o25: y = {a[20:0], a[31:21]};
			5'o26: y = {a[21:0], a[31:22]};
			5'o27: y = {a[22:0], a[31:23]};
			5'o30: y = {a[23:0], a[31:24]};
			5'o31: y = {a[24:0], a[31:25]};
			5'o32: y = {a[25:0], a[31:26]};
			5'o33: y = {a[26:0], a[31:27]};
			5'o34: y = {a[27:0], a[31:28]};
			5'o35: y = {a[28:0], a[31:29]};
			5'o36: y = {a[29:0], a[31:30]};
			5'o37: y = {a[30:0], a[31]};
			default: y = a;
		endcase
	  else
		  case(amt)//right
			5'o0: y = a;
			5'o37: y = {a[0], a[31:1]};
			5'o36: y = {a[1:0], a[31:2]};
			5'o35: y = {a[2:0], a[31:3]};
			5'o34: y = {a[3:0], a[31:4]};
			5'o33: y = {a[4:0], a[31:5]};
			5'o32: y = {a[5:0], a[31:6]};
			5'o31: y = {a[6:0], a[31:7]};
			5'o30: y = {a[7:0], a[31:8]};
			5'o27: y = {a[8:0], a[31:9]};
			5'o26: y = {a[9:0], a[31:10]};
			5'o25: y = {a[10:0], a[31:11]};
			5'o24: y = {a[11:0], a[31:12]};
			5'o23: y = {a[12:0], a[31:13]};
			5'o22: y = {a[13:0], a[31:14]};
			5'o21: y = {a[14:0], a[31:15]};
			5'o20: y = {a[15:0], a[31:16]};
			5'o17: y = {a[16:0], a[31:17]};
			5'o16: y = {a[17:0], a[31:18]};
			5'o15: y = {a[18:0], a[31:19]};
			5'o14: y = {a[19:0], a[31:20]};
			5'o13: y = {a[20:0], a[31:21]};
			5'o12: y = {a[21:0], a[31:22]};
			5'o11: y = {a[22:0], a[31:23]};
			5'o10: y = {a[23:0], a[31:24]};
			5'o7: y = {a[24:0], a[31:25]};
			5'o6: y = {a[25:0], a[31:26]};
			5'o5: y = {a[26:0], a[31:27]};
			5'o4: y = {a[27:0], a[31:28]};
			5'o3: y = {a[28:0], a[31:29]};
			5'o2: y = {a[29:0], a[31:30]};
			5'o1: y = {a[30:0], a[31]};
			default: y = a;
			endcase
  end
endmodule
